module instructionmemory (
	output reg [31:0] saida,
	input Clk,
	input [9:0] endereco
);	
	
	reg [31:0] memoria [0:1023];
		
	integer i;
	
	always @(posedge Clk) begin
		saida <= memoria[endereco];
	end

/*	
#define A 0x1500
#define B 0x1501
#define C 0x1502
#define D 0x1503
#define END 0x18FF

lw $r0, A(r31)
lw $r1, B(r31)
lw $r2, C(r31)
lw $r3, D(r31)

mul $r4, $r0, $r1
add $r5, $r2, $r3
sub $r6, $r4, $r5

sw $r6, END(r31)


Traduzindo para instruções em binário:

001000_11111_00000_0001-0101-0000-0000
001000_11111_00001_0001-0101-0000-0001
001000_11111_00010_0001-0101-0000-0010
001000_11111_00011_0001-0101-0000-0011

000111_00000_00001_00100_01010_110010
000111_00010_00011_00101_01010_100000
000111_00100_00101_00110_01010_100010

001001_11111_00110_0001-1000-1111-1111



Bolhas:

and r30, r30, r30
or r29, r29, r29

000111_11110_11110_11110_01010_100100
000111_11101_11101_11101_01010_100101
*/
	
	initial begin
		memoria[0]=32'b001000_11111_00000_0001010100000000;
		memoria[1]=32'b001000_11111_00001_0001010100000001;
		memoria[2]=32'b001000_11111_00010_0001010100000010;
		memoria[3]=32'b001000_11111_00011_0001010100000011;
		
		memoria[4]=32'b000111_00000_00001_00100_01010_110010;
		memoria[5]=32'b000111_00010_00011_00101_01010_100000;
		memoria[6]=32'b000111_00100_00101_00110_01010_100010;

		memoria[7]=32'b001001_11111_00110_0001100011111111;
		
		//Mesmo programa mas com bolhas:
		memoria[8]=32'b001000_11111_00000_0001010100000000;
		memoria[9]=32'b001000_11111_00001_0001010100000001;
		memoria[10]=32'b001000_11111_00010_0001010100000010;
		memoria[11]=32'b001000_11111_00011_0001010100000011;
		
		memoria[12]=32'b000111_00000_00001_00100_01010_110010;
		memoria[13]=32'b000111_00010_00011_00101_01010_100000;
		memoria[14]=32'b000111_11110_11110_11110_01010_100100;//bolhaAnd
		memoria[15]=32'b000111_11110_11110_11110_01010_100100;//bolhaAnd
		memoria[16]=32'b000111_11110_11110_11110_01010_100100;//bolhaAnd
		memoria[17]=32'b000111_00100_00101_00110_01010_100010;
		
		memoria[18]=32'b000111_11101_11101_11101_01010_100101;//bolhaOr
		memoria[19]=32'b000111_11101_11101_11101_01010_100101;//bolhaOr
		memoria[20]=32'b000111_11101_11101_11101_01010_100101;//bolhaOr
		memoria[21]=32'b001001_11111_00110_0001100011111111;
	
		for(i = 22; i < 1024;i = i+1) 
			memoria[i] = 32'b0;
	end

endmodule 

