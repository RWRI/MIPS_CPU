module pll();
endmodule
